
module ISSP (
	probe,
	source_clk,
	source);	

	input	[61:0]	probe;
	input		source_clk;
	output	[92:0]	source;
endmodule
