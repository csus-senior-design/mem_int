
module ISSP (
	source,
	probe,
	source_clk);	

	output	[1:0]	source;
	input	[6:0]	probe;
	input		source_clk;
endmodule
